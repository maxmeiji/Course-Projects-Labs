module labsix3(LEDR,SW,KEY,CLOCK_50,HEX0,HEX1,HEX2,HEX3);
	input [3:0]KEY;
	output reg [0:0] LEDR;
	input CLOCK_50;
	output [6:0]HEX0;
	output [6:0]HEX1;
	output [6:0]HEX2;
	output [6:0]HEX3;
	reg [30:0]Q,D;
	reg [3:0]s,start,sig,sig2,R4,R3,R2,R1;
	input [9:0]SW;
	
	
	always @(posedge CLOCK_50)begin
	if(start==1)begin
		if(Q == s*50000000)begin
			Q <= 0;
			sig<=1;
			LEDR[0]<=1;
		
		end
		else begin
		Q<=Q+1;
	
		end
			
		end
	if(start==0) begin
		LEDR[0]<=0;
		sig<=0;
	end
	
	if(sig==1)begin
		
		if(D == 50000)begin
			D <= 0;
			if(R1==9) begin
				R1<=0;
				if(R2==9) begin
					R2<=0;
					if(R3==9) begin
						R3<=0;
						R4<=R4+1;
					end
					
					else begin
						R3<=R3+1;
					end
				end
				else begin
					R2<=R2+1;
				end
			end
			
			else begin
				R1<=R1+1;
			end
			end
		else begin
			D<=D+1;
		end
			end
	if(sig==0 && sig2==0) begin	
				R1<=0;
				R2<=0;
				R3<=0;
				R4<=0;
			end
			
			
			
		end


	always@(negedge KEY[0], negedge KEY[3]) begin
		if(KEY[0]==0) begin
			start<=1;
			s<=SW[3:0];
			sig2=0;
		end
		if(KEY[3]==0) begin
			start<=0;
			sig2<=1;
		end
	end

	hexto7segment s2(R4,HEX3);
	hexto7segment s3(R3,HEX2);
	hexto7segment s4(R2,HEX1);
	hexto7segment s5(R1,HEX0);

	endmodule

module hexto7segment (
   input [3:0] iDIG,
   output reg [6:0] oSEG
	 );
 
 always@(iDIG) begin
   case(iDIG)
     4'b0001: oSEG = 7'b1111001;
	  4'b0010: oSEG = 7'b0100100;  // ---t----     4'h2: oSEG = 7'b0100100;  // |      |
     4'b0011: oSEG = 7'b0110000;  // lt    rt
     4'b0100: oSEG = 7'b0011001;  // |      |
     4'b0101: oSEG = 7'b0010010;  // ---m----
     4'b0110: oSEG = 7'b0000010;  // |      |
     4'b0111: oSEG = 7'b1111000;  // lb    rb
     4'b1000: oSEG = 7'b0000000;  // |      |
     4'b1001: oSEG = 7'b0011000;  // ---b----
     4'b0000: oSEG = 7'b1000000;
   endcase
 end
 
endmodule